`define IDLE_MODE 0
`define FC_MODE 1
`define CONV_MODE 2
`define EMPTY_MODE 3
