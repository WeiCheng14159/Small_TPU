// This file include all user-defined package

`include "accelerator_pkg.sv"
`include "systolic_array_pkg.sv"
`include "single_port_ram_pkg.sv"
